Usage: scripts/generate_image_rom.py <input_png> <output_file>
